//module Table_FSM(
//	
//);
//
//endmodule
module Memory_Controller ()

endmodule
